program mem_program();
  mem_env env;
 initial begin
    env=new();
    env.run();
end

endprogram
