
`include "memory.v"
`include "mem_common.sv"
`include "mem_intf.sv"
`include "mem_assert.sv"
`include "mem_tx.sv"
`include "mem_gen.sv"
`include "mem_bfm.sv"
`include "mem_cov.sv"
`include "mem_mon.sv"
`include "mem_sbd.sv"
`include "mem_agt.sv"
`include "mem_env.sv"
//`include "mem_program.sv"
`include "mem_top.sv"

//https://edaplayground.com/x/MWqp

//0https://edaplayground.com/x/ZrMP

